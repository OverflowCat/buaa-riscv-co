module control(
);


endmodule


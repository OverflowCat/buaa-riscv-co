module control(
       input[31:0] instr,
       output      branch,
       output      memread,
       output      memtoreg,
       output[3:0] aluctrl,
       output      alusrc,
       output      memwrite,
       output      regwrite 
);

//请在这里补充你的控制器代码

endmodule


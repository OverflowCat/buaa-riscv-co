module data_path (

);


endmodule //data_path
















module data_ram(
    input clk,
    input WE,
    input RE,
    input[31:0] A,
    input[31:0] WD,
    output[31:0] RD
);

//请在这里补充你的数据存储器代码

endmodule

module imm_gen(
    input [31:0] instr,
    output[31:0] imm
);

//请在这里补充你的立即数生成模块代码

endmodule

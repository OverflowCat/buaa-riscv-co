module alu (
    input  wire [32-1:0] A,
    input  wire [32-1:0] B,
    input  wire [4-1 :0] ALUCtrl,
    output wire          ZERO,
    output wire [32-1:0] Y
);

//请在这里补充你的ALU实现代码

endmodule
module regfile (
);


reg[32-1:0]   rf[32-1:0];


endmodule //regfile


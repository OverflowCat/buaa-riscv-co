module pc_rom(
);

reg[32-1:0] cpu_instr_rom[2047:0];


endmodule

module alu (
);


endmodule //alu
module data_ram(
    
);


endmodule

module core_top(
             
    input  wire  clk,
    input  wire  rst_n
);

data_path u_data_path (
     
);

control  u_controller(
       
);

endmodule

module regfile (
    input  wire         clk,
    input  wire         WE,
    input  wire[5-1:0]  A1,
    input  wire[5-1:0]  A2,
    input  wire[5-1:0]  A3,
    input  wire[32-1:0] WD3,
    output wire[32-1:0] RD1,
    output wire[32-1:0] RD2
);

//请在这里补充你设计的寄存器堆代码

endmodule

